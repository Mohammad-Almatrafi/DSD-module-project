module FSM_Rx (
    clk,
    rst_n,
    count15_rst_n,
    count15_en,
    count_size_rst_n,
    count_size_en,
    shift_reg_en,
    shift_reg_rst_n
);
  input clk, rst_n;
  output count15_en, count15_rst_n, count_size_en, count_size_rst_n, shift_reg_en, shift_reg_rst_n;





endmodule
