module Datapath_Rx (
    clk,
    rst_n,
    counter_sample_rst_n,
    counter_sample_en,
    counter_size_en,
    counter_size_rst_n,


);

  // shift reg is needed

endmodule
