module Datapath_Rx ();




endmodule
